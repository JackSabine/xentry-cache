`include "dcache_test.sv"
