module no_test();

initial begin
  $finish();
end

endmodule
