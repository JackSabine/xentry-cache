`include "dcache_load_test.sv"
`include "dcache_load_hit_test.sv"
`include "dcache_clflush_test.sv"
