typedef uvm_sequencer #(reset_transaction) reset_sequencer;
