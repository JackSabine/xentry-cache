`include "dcache_load_test.sv"
`include "dcache_load_hit_test.sv"
`include "dcache_clflush_test.sv"
`include "dcache_store_test.sv"
`include "dcache_full_test.sv"
`include "icache_full_test.sv"
