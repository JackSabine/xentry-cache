typedef uvm_sequencer #(memory_transaction) memory_sequencer;