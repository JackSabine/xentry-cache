`include "memory_simple_test.sv"
