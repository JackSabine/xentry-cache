`include "icache_basic_test.sv"
