`include "cache_base_test.sv"
`include "icache_basic_test.sv"
