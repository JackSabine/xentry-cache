`ifndef MACROS__SVH
  `define MACROS__SVH

`define WORD        (32)
`define HALF        (16)
`define BYTE        (8)
`define REG_BITS    (5)
`define NUM_REGS    (32)

typedef int unsigned uint32_t;

`endif