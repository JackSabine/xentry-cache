`include "dcache_load_test.sv"
`include "dcache_store_test.sv"
