import "DPI-C" function string get_environment_variable(string env_name);
