typedef uvm_sequencer #(memory_transaction) cache_req_sequencer;
